----------------------------------------------------------------------------------
--                                 _             _
--                                | |_  ___ _ __(_)__ _
--                                | ' \/ -_) '_ \ / _` |
--                                |_||_\___| .__/_\__,_|
--                                         |_|
--
----------------------------------------------------------------------------------
--
-- Company: hepia
-- Author: Orphee Antoniadis <orphee.antoniadis@hesge.ch>
--
-- Module Name: tb_zybo_pcam5c_zynqps - arch
-- Target Device: digilentinc.com:zybo-z7-20:part0:1.0 xc7z020clg400-1
-- Tool version: 2020.2
-- Description: Testbench for zybo_pcam5c_zynqps
--
-- Last update: 2021-08-10 12:21:11
--
---------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_zybo_pcam5c_zynqps is
end tb_zybo_pcam5c_zynqps;


architecture behavioral of tb_zybo_pcam5c_zynqps is

begin

end behavioral;
